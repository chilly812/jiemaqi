module ycc_rgb_convert (dataa,
		 datab,
                 result                      	
		);

input [31:0] dataa ; // 32 bit write data line
input [31:0] datab ; // 32 bit write data line
output reg [31:0] result ;

reg [31:0] dataa_reg ;
reg [31:0] datab_reg ;

reg [7:0] y;
reg [7:0] cr;
reg [7:0] cb;

reg [7:0] R;
reg [7:0] G;
reg [7:0] B;

reg signed [31:0] cr_r [255:0];
reg signed [31:0] cr_g [255:0];
reg signed [31:0] cb_b [255:0];
reg signed [31:0] cb_g [255:0];


initial begin

cr_r[0] = -32'sd179;
cr_r[1] = -32'sd178;
cr_r[2] = -32'sd177;
cr_r[3] = -32'sd175;
cr_r[4] = -32'sd174;
cr_r[5] = -32'sd172;
cr_r[6] = -32'sd171;
cr_r[7] = -32'sd170;
cr_r[8] = -32'sd168;
cr_r[9] = -32'sd167;
cr_r[10] = -32'sd165;
cr_r[11] = -32'sd164;
cr_r[12] = -32'sd163;
cr_r[13] = -32'sd161;
cr_r[14] = -32'sd160;
cr_r[15] = -32'sd158;
cr_r[16] = -32'sd157;
cr_r[17] = -32'sd156;
cr_r[18] = -32'sd154;
cr_r[19] = -32'sd153;
cr_r[20] = -32'sd151;
cr_r[21] = -32'sd150;
cr_r[22] = -32'sd149;
cr_r[23] = -32'sd147;
cr_r[24] = -32'sd146;
cr_r[25] = -32'sd144;
cr_r[26] = -32'sd143;
cr_r[27] = -32'sd142;
cr_r[28] = -32'sd140;
cr_r[29] = -32'sd139;
cr_r[30] = -32'sd137;
cr_r[31] = -32'sd136;
cr_r[32] = -32'sd135;
cr_r[33] = -32'sd133;
cr_r[34] = -32'sd132;
cr_r[35] = -32'sd130;
cr_r[36] = -32'sd129;
cr_r[37] = -32'sd128;
cr_r[38] = -32'sd126;
cr_r[39] = -32'sd125;
cr_r[40] = -32'sd123;
cr_r[41] = -32'sd122;
cr_r[42] = -32'sd121;
cr_r[43] = -32'sd119;
cr_r[44] = -32'sd118;
cr_r[45] = -32'sd116;
cr_r[46] = -32'sd115;
cr_r[47] = -32'sd114;
cr_r[48] = -32'sd112;
cr_r[49] = -32'sd111;
cr_r[50] = -32'sd109;
cr_r[51] = -32'sd108;
cr_r[52] = -32'sd107;
cr_r[53] = -32'sd105;
cr_r[54] = -32'sd104;
cr_r[55] = -32'sd102;
cr_r[56] = -32'sd101;
cr_r[57] = -32'sd100;
cr_r[58] = -32'sd98;
cr_r[59] = -32'sd97;
cr_r[60] = -32'sd95;
cr_r[61] = -32'sd94;
cr_r[62] = -32'sd93;
cr_r[63] = -32'sd91;
cr_r[64] = -32'sd90;
cr_r[65] = -32'sd88;
cr_r[66] = -32'sd87;
cr_r[67] = -32'sd86;
cr_r[68] = -32'sd84;
cr_r[69] = -32'sd83;
cr_r[70] = -32'sd81;
cr_r[71] = -32'sd80;
cr_r[72] = -32'sd79;
cr_r[73] = -32'sd77;
cr_r[74] = -32'sd76;
cr_r[75] = -32'sd74;
cr_r[76] = -32'sd73;
cr_r[77] = -32'sd72;
cr_r[78] = -32'sd70;
cr_r[79] = -32'sd69;
cr_r[80] = -32'sd67;
cr_r[81] = -32'sd66;
cr_r[82] = -32'sd64;
cr_r[83] = -32'sd63;
cr_r[84] = -32'sd62;
cr_r[85] = -32'sd60;
cr_r[86] = -32'sd59;
cr_r[87] = -32'sd57;
cr_r[88] = -32'sd56;
cr_r[89] = -32'sd55;
cr_r[90] = -32'sd53;
cr_r[91] = -32'sd52;
cr_r[92] = -32'sd50;
cr_r[93] = -32'sd49;
cr_r[94] = -32'sd48;
cr_r[95] = -32'sd46;
cr_r[96] = -32'sd45;
cr_r[97] = -32'sd43;
cr_r[98] = -32'sd42;
cr_r[99] = -32'sd41;
cr_r[100] = -32'sd39;
cr_r[101] = -32'sd38;
cr_r[102] = -32'sd36;
cr_r[103] = -32'sd35;
cr_r[104] = -32'sd34;
cr_r[105] = -32'sd32;
cr_r[106] = -32'sd31;
cr_r[107] = -32'sd29;
cr_r[108] = -32'sd28;
cr_r[109] = -32'sd27;
cr_r[110] = -32'sd25;
cr_r[111] = -32'sd24;
cr_r[112] = -32'sd22;
cr_r[113] = -32'sd21;
cr_r[114] = -32'sd20;
cr_r[115] = -32'sd18;
cr_r[116] = -32'sd17;
cr_r[117] = -32'sd15;
cr_r[118] = -32'sd14;
cr_r[119] = -32'sd13;
cr_r[120] = -32'sd11;
cr_r[121] = -32'sd10;
cr_r[122] = -32'sd8;
cr_r[123] = -32'sd7;
cr_r[124] = -32'sd6;
cr_r[125] = -32'sd4;
cr_r[126] = -32'sd3;
cr_r[127] = -32'sd1;
cr_r[128] = -32'sd0;
cr_r[129] = 32'sd1;
cr_r[130] = 32'sd3;
cr_r[131] = 32'sd4;
cr_r[132] = 32'sd6;
cr_r[133] = 32'sd7;
cr_r[134] = 32'sd8;
cr_r[135] = 32'sd10;
cr_r[136] = 32'sd11;
cr_r[137] = 32'sd13;
cr_r[138] = 32'sd14;
cr_r[139] = 32'sd15;
cr_r[140] = 32'sd17;
cr_r[141] = 32'sd18;
cr_r[142] = 32'sd20;
cr_r[143] = 32'sd21;
cr_r[144] = 32'sd22;
cr_r[145] = 32'sd24;
cr_r[146] = 32'sd25;
cr_r[147] = 32'sd27;
cr_r[148] = 32'sd28;
cr_r[149] = 32'sd29;
cr_r[150] = 32'sd31;
cr_r[151] = 32'sd32;
cr_r[152] = 32'sd34;
cr_r[153] = 32'sd35;
cr_r[154] = 32'sd36;
cr_r[155] = 32'sd38;
cr_r[156] = 32'sd39;
cr_r[157] = 32'sd41;
cr_r[158] = 32'sd42;
cr_r[159] = 32'sd43;
cr_r[160] = 32'sd45;
cr_r[161] = 32'sd46;
cr_r[162] = 32'sd48;
cr_r[163] = 32'sd49;
cr_r[164] = 32'sd50;
cr_r[165] = 32'sd52;
cr_r[166] = 32'sd53;
cr_r[167] = 32'sd55;
cr_r[168] = 32'sd56;
cr_r[169] = 32'sd57;
cr_r[170] = 32'sd59;
cr_r[171] = 32'sd60;
cr_r[172] = 32'sd62;
cr_r[173] = 32'sd63;
cr_r[174] = 32'sd64;
cr_r[175] = 32'sd66;
cr_r[176] = 32'sd67;
cr_r[177] = 32'sd69;
cr_r[178] = 32'sd70;
cr_r[179] = 32'sd72;
cr_r[180] = 32'sd73;
cr_r[181] = 32'sd74;
cr_r[182] = 32'sd76;
cr_r[183] = 32'sd77;
cr_r[184] = 32'sd79;
cr_r[185] = 32'sd80;
cr_r[186] = 32'sd81;
cr_r[187] = 32'sd83;
cr_r[188] = 32'sd84;
cr_r[189] = 32'sd86;
cr_r[190] = 32'sd87;
cr_r[191] = 32'sd88;
cr_r[192] = 32'sd90;
cr_r[193] = 32'sd91;
cr_r[194] = 32'sd93;
cr_r[195] = 32'sd94;
cr_r[196] = 32'sd95;
cr_r[197] = 32'sd97;
cr_r[198] = 32'sd98;
cr_r[199] = 32'sd100;
cr_r[200] = 32'sd101;
cr_r[201] = 32'sd102;
cr_r[202] = 32'sd104;
cr_r[203] = 32'sd105;
cr_r[204] = 32'sd107;
cr_r[205] = 32'sd108;
cr_r[206] = 32'sd109;
cr_r[207] = 32'sd111;
cr_r[208] = 32'sd112;
cr_r[209] = 32'sd114;
cr_r[210] = 32'sd115;
cr_r[211] = 32'sd116;
cr_r[212] = 32'sd118;
cr_r[213] = 32'sd119;
cr_r[214] = 32'sd121;
cr_r[215] = 32'sd122;
cr_r[216] = 32'sd123;
cr_r[217] = 32'sd125;
cr_r[218] = 32'sd126;
cr_r[219] = 32'sd128;
cr_r[220] = 32'sd129;
cr_r[221] = 32'sd130;
cr_r[222] = 32'sd132;
cr_r[223] = 32'sd133;
cr_r[224] = 32'sd135;
cr_r[225] = 32'sd136;
cr_r[226] = 32'sd137;
cr_r[227] = 32'sd139;
cr_r[228] = 32'sd140;
cr_r[229] = 32'sd142;
cr_r[230] = 32'sd143;
cr_r[231] = 32'sd144;
cr_r[232] = 32'sd146;
cr_r[233] = 32'sd147;
cr_r[234] = 32'sd149;
cr_r[235] = 32'sd150;
cr_r[236] = 32'sd151;
cr_r[237] = 32'sd153;
cr_r[238] = 32'sd154;
cr_r[239] = 32'sd156;
cr_r[240] = 32'sd157;
cr_r[241] = 32'sd158;
cr_r[242] = 32'sd160;
cr_r[243] = 32'sd161;
cr_r[244] = 32'sd163;
cr_r[245] = 32'sd164;
cr_r[246] = 32'sd165;
cr_r[247] = 32'sd167;
cr_r[248] = 32'sd168;
cr_r[249] = 32'sd170;
cr_r[250] = 32'sd171;
cr_r[251] = 32'sd172;
cr_r[252] = 32'sd174;
cr_r[253] = 32'sd175;
cr_r[254] = 32'sd177;
cr_r[255] = 32'sd178;


cr_g[0] = 32'sd5990656;
cr_g[1] = 32'sd5943854;
cr_g[2] = 32'sd5897052;
cr_g[3] = 32'sd5850250;
cr_g[4] = 32'sd5803448;
cr_g[5] = 32'sd5756646;
cr_g[6] = 32'sd5709844;
cr_g[7] = 32'sd5663042;
cr_g[8] = 32'sd5616240;
cr_g[9] = 32'sd5569438;
cr_g[10] = 32'sd5522636;
cr_g[11] = 32'sd5475834;
cr_g[12] = 32'sd5429032;
cr_g[13] = 32'sd5382230;
cr_g[14] = 32'sd5335428;
cr_g[15] = 32'sd5288626;
cr_g[16] = 32'sd5241824;
cr_g[17] = 32'sd5195022;
cr_g[18] = 32'sd5148220;
cr_g[19] = 32'sd5101418;
cr_g[20] = 32'sd5054616;
cr_g[21] = 32'sd5007814;
cr_g[22] = 32'sd4961012;
cr_g[23] = 32'sd4914210;
cr_g[24] = 32'sd4867408;
cr_g[25] = 32'sd4820606;
cr_g[26] = 32'sd4773804;
cr_g[27] = 32'sd4727002;
cr_g[28] = 32'sd4680200;
cr_g[29] = 32'sd4633398;
cr_g[30] = 32'sd4586596;
cr_g[31] = 32'sd4539794;
cr_g[32] = 32'sd4492992;
cr_g[33] = 32'sd4446190;
cr_g[34] = 32'sd4399388;
cr_g[35] = 32'sd4352586;
cr_g[36] = 32'sd4305784;
cr_g[37] = 32'sd4258982;
cr_g[38] = 32'sd4212180;
cr_g[39] = 32'sd4165378;
cr_g[40] = 32'sd4118576;
cr_g[41] = 32'sd4071774;
cr_g[42] = 32'sd4024972;
cr_g[43] = 32'sd3978170;
cr_g[44] = 32'sd3931368;
cr_g[45] = 32'sd3884566;
cr_g[46] = 32'sd3837764;
cr_g[47] = 32'sd3790962;
cr_g[48] = 32'sd3744160;
cr_g[49] = 32'sd3697358;
cr_g[50] = 32'sd3650556;
cr_g[51] = 32'sd3603754;
cr_g[52] = 32'sd3556952;
cr_g[53] = 32'sd3510150;
cr_g[54] = 32'sd3463348;
cr_g[55] = 32'sd3416546;
cr_g[56] = 32'sd3369744;
cr_g[57] = 32'sd3322942;
cr_g[58] = 32'sd3276140;
cr_g[59] = 32'sd3229338;
cr_g[60] = 32'sd3182536;
cr_g[61] = 32'sd3135734;
cr_g[62] = 32'sd3088932;
cr_g[63] = 32'sd3042130;
cr_g[64] = 32'sd2995328;
cr_g[65] = 32'sd2948526;
cr_g[66] = 32'sd2901724;
cr_g[67] = 32'sd2854922;
cr_g[68] = 32'sd2808120;
cr_g[69] = 32'sd2761318;
cr_g[70] = 32'sd2714516;
cr_g[71] = 32'sd2667714;
cr_g[72] = 32'sd2620912;
cr_g[73] = 32'sd2574110;
cr_g[74] = 32'sd2527308;
cr_g[75] = 32'sd2480506;
cr_g[76] = 32'sd2433704;
cr_g[77] = 32'sd2386902;
cr_g[78] = 32'sd2340100;
cr_g[79] = 32'sd2293298;
cr_g[80] = 32'sd2246496;
cr_g[81] = 32'sd2199694;
cr_g[82] = 32'sd2152892;
cr_g[83] = 32'sd2106090;
cr_g[84] = 32'sd2059288;
cr_g[85] = 32'sd2012486;
cr_g[86] = 32'sd1965684;
cr_g[87] = 32'sd1918882;
cr_g[88] = 32'sd1872080;
cr_g[89] = 32'sd1825278;
cr_g[90] = 32'sd1778476;
cr_g[91] = 32'sd1731674;
cr_g[92] = 32'sd1684872;
cr_g[93] = 32'sd1638070;
cr_g[94] = 32'sd1591268;
cr_g[95] = 32'sd1544466;
cr_g[96] = 32'sd1497664;
cr_g[97] = 32'sd1450862;
cr_g[98] = 32'sd1404060;
cr_g[99] = 32'sd1357258;
cr_g[100] = 32'sd1310456;
cr_g[101] = 32'sd1263654;
cr_g[102] = 32'sd1216852;
cr_g[103] = 32'sd1170050;
cr_g[104] = 32'sd1123248;
cr_g[105] = 32'sd1076446;
cr_g[106] = 32'sd1029644;
cr_g[107] = 32'sd982842;
cr_g[108] = 32'sd936040;
cr_g[109] = 32'sd889238;
cr_g[110] = 32'sd842436;
cr_g[111] = 32'sd795634;
cr_g[112] = 32'sd748832;
cr_g[113] = 32'sd702030;
cr_g[114] = 32'sd655228;
cr_g[115] = 32'sd608426;
cr_g[116] = 32'sd561624;
cr_g[117] = 32'sd514822;
cr_g[118] = 32'sd468020;
cr_g[119] = 32'sd421218;
cr_g[120] = 32'sd374416;
cr_g[121] = 32'sd327614;
cr_g[122] = 32'sd280812;
cr_g[123] = 32'sd234010;
cr_g[124] = 32'sd187208;
cr_g[125] = 32'sd140406;
cr_g[126] = 32'sd93604;
cr_g[127] = 32'sd46802;
cr_g[128] = 32'sd0;
cr_g[129] = -32'sd46802;
cr_g[130] = -32'sd93604;
cr_g[131] = -32'sd140406;
cr_g[132] = -32'sd187208;
cr_g[133] = -32'sd234010;
cr_g[134] = -32'sd280812;
cr_g[135] = -32'sd327614;
cr_g[136] = -32'sd374416;
cr_g[137] = -32'sd421218;
cr_g[138] = -32'sd468020;
cr_g[139] = -32'sd514822;
cr_g[140] = -32'sd561624;
cr_g[141] = -32'sd608426;
cr_g[142] = -32'sd655228;
cr_g[143] = -32'sd702030;
cr_g[144] = -32'sd748832;
cr_g[145] = -32'sd795634;
cr_g[146] = -32'sd842436;
cr_g[147] = -32'sd889238;
cr_g[148] = -32'sd936040;
cr_g[149] = -32'sd982842;
cr_g[150] = -32'sd1029644;
cr_g[151] = -32'sd1076446;
cr_g[152] = -32'sd1123248;
cr_g[153] = -32'sd1170050;
cr_g[154] = -32'sd1216852;
cr_g[155] = -32'sd1263654;
cr_g[156] = -32'sd1310456;
cr_g[157] = -32'sd1357258;
cr_g[158] = -32'sd1404060;
cr_g[159] = -32'sd1450862;
cr_g[160] = -32'sd1497664;
cr_g[161] = -32'sd1544466;
cr_g[162] = -32'sd1591268;
cr_g[163] = -32'sd1638070;
cr_g[164] = -32'sd1684872;
cr_g[165] = -32'sd1731674;
cr_g[166] = -32'sd1778476;
cr_g[167] = -32'sd1825278;
cr_g[168] = -32'sd1872080;
cr_g[169] = -32'sd1918882;
cr_g[170] = -32'sd1965684;
cr_g[171] = -32'sd2012486;
cr_g[172] = -32'sd2059288;
cr_g[173] = -32'sd2106090;
cr_g[174] = -32'sd2152892;
cr_g[175] = -32'sd2199694;
cr_g[176] = -32'sd2246496;
cr_g[177] = -32'sd2293298;
cr_g[178] = -32'sd2340100;
cr_g[179] = -32'sd2386902;
cr_g[180] = -32'sd2433704;
cr_g[181] = -32'sd2480506;
cr_g[182] = -32'sd2527308;
cr_g[183] = -32'sd2574110;
cr_g[184] = -32'sd2620912;
cr_g[185] = -32'sd2667714;
cr_g[186] = -32'sd2714516;
cr_g[187] = -32'sd2761318;
cr_g[188] = -32'sd2808120;
cr_g[189] = -32'sd2854922;
cr_g[190] = -32'sd2901724;
cr_g[191] = -32'sd2948526;
cr_g[192] = -32'sd2995328;
cr_g[193] = -32'sd3042130;
cr_g[194] = -32'sd3088932;
cr_g[195] = -32'sd3135734;
cr_g[196] = -32'sd3182536;
cr_g[197] = -32'sd3229338;
cr_g[198] = -32'sd3276140;
cr_g[199] = -32'sd3322942;
cr_g[200] = -32'sd3369744;
cr_g[201] = -32'sd3416546;
cr_g[202] = -32'sd3463348;
cr_g[203] = -32'sd3510150;
cr_g[204] = -32'sd3556952;
cr_g[205] = -32'sd3603754;
cr_g[206] = -32'sd3650556;
cr_g[207] = -32'sd3697358;
cr_g[208] = -32'sd3744160;
cr_g[209] = -32'sd3790962;
cr_g[210] = -32'sd3837764;
cr_g[211] = -32'sd3884566;
cr_g[212] = -32'sd3931368;
cr_g[213] = -32'sd3978170;
cr_g[214] = -32'sd4024972;
cr_g[215] = -32'sd4071774;
cr_g[216] = -32'sd4118576;
cr_g[217] = -32'sd4165378;
cr_g[218] = -32'sd4212180;
cr_g[219] = -32'sd4258982;
cr_g[220] = -32'sd4305784;
cr_g[221] = -32'sd4352586;
cr_g[222] = -32'sd4399388;
cr_g[223] = -32'sd4446190;
cr_g[224] = -32'sd4492992;
cr_g[225] = -32'sd4539794;
cr_g[226] = -32'sd4586596;
cr_g[227] = -32'sd4633398;
cr_g[228] = -32'sd4680200;
cr_g[229] = -32'sd4727002;
cr_g[230] = -32'sd4773804;
cr_g[231] = -32'sd4820606;
cr_g[232] = -32'sd4867408;
cr_g[233] = -32'sd4914210;
cr_g[234] = -32'sd4961012;
cr_g[235] = -32'sd5007814;
cr_g[236] = -32'sd5054616;
cr_g[237] = -32'sd5101418;
cr_g[238] = -32'sd5148220;
cr_g[239] = -32'sd5195022;
cr_g[240] = -32'sd5241824;
cr_g[241] = -32'sd5288626;
cr_g[242] = -32'sd5335428;
cr_g[243] = -32'sd5382230;
cr_g[244] = -32'sd5429032;
cr_g[245] = -32'sd5475834;
cr_g[246] = -32'sd5522636;
cr_g[247] = -32'sd5569438;
cr_g[248] = -32'sd5616240;
cr_g[249] = -32'sd5663042;
cr_g[250] = -32'sd5709844;
cr_g[251] = -32'sd5756646;
cr_g[252] = -32'sd5803448;
cr_g[253] = -32'sd5850250;
cr_g[254] = -32'sd5897052;
cr_g[255] = -32'sd5943854;


cb_b[0] = -32'sd227;
cb_b[1] = -32'sd225;
cb_b[2] = -32'sd223;
cb_b[3] = -32'sd222;
cb_b[4] = -32'sd220;
cb_b[5] = -32'sd218;
cb_b[6] = -32'sd216;
cb_b[7] = -32'sd214;
cb_b[8] = -32'sd213;
cb_b[9] = -32'sd211;
cb_b[10] = -32'sd209;
cb_b[11] = -32'sd207;
cb_b[12] = -32'sd206;
cb_b[13] = -32'sd204;
cb_b[14] = -32'sd202;
cb_b[15] = -32'sd200;
cb_b[16] = -32'sd198;
cb_b[17] = -32'sd197;
cb_b[18] = -32'sd195;
cb_b[19] = -32'sd193;
cb_b[20] = -32'sd191;
cb_b[21] = -32'sd190;
cb_b[22] = -32'sd188;
cb_b[23] = -32'sd186;
cb_b[24] = -32'sd184;
cb_b[25] = -32'sd183;
cb_b[26] = -32'sd181;
cb_b[27] = -32'sd179;
cb_b[28] = -32'sd177;
cb_b[29] = -32'sd175;
cb_b[30] = -32'sd174;
cb_b[31] = -32'sd172;
cb_b[32] = -32'sd170;
cb_b[33] = -32'sd168;
cb_b[34] = -32'sd167;
cb_b[35] = -32'sd165;
cb_b[36] = -32'sd163;
cb_b[37] = -32'sd161;
cb_b[38] = -32'sd159;
cb_b[39] = -32'sd158;
cb_b[40] = -32'sd156;
cb_b[41] = -32'sd154;
cb_b[42] = -32'sd152;
cb_b[43] = -32'sd151;
cb_b[44] = -32'sd149;
cb_b[45] = -32'sd147;
cb_b[46] = -32'sd145;
cb_b[47] = -32'sd144;
cb_b[48] = -32'sd142;
cb_b[49] = -32'sd140;
cb_b[50] = -32'sd138;
cb_b[51] = -32'sd136;
cb_b[52] = -32'sd135;
cb_b[53] = -32'sd133;
cb_b[54] = -32'sd131;
cb_b[55] = -32'sd129;
cb_b[56] = -32'sd128;
cb_b[57] = -32'sd126;
cb_b[58] = -32'sd124;
cb_b[59] = -32'sd122;
cb_b[60] = -32'sd120;
cb_b[61] = -32'sd119;
cb_b[62] = -32'sd117;
cb_b[63] = -32'sd115;
cb_b[64] = -32'sd113;
cb_b[65] = -32'sd112;
cb_b[66] = -32'sd110;
cb_b[67] = -32'sd108;
cb_b[68] = -32'sd106;
cb_b[69] = -32'sd105;
cb_b[70] = -32'sd103;
cb_b[71] = -32'sd101;
cb_b[72] = -32'sd99;
cb_b[73] = -32'sd97;
cb_b[74] = -32'sd96;
cb_b[75] = -32'sd94;
cb_b[76] = -32'sd92;
cb_b[77] = -32'sd90;
cb_b[78] = -32'sd89;
cb_b[79] = -32'sd87;
cb_b[80] = -32'sd85;
cb_b[81] = -32'sd83;
cb_b[82] = -32'sd82;
cb_b[83] = -32'sd80;
cb_b[84] = -32'sd78;
cb_b[85] = -32'sd76;
cb_b[86] = -32'sd74;
cb_b[87] = -32'sd73;
cb_b[88] = -32'sd71;
cb_b[89] = -32'sd69;
cb_b[90] = -32'sd67;
cb_b[91] = -32'sd66;
cb_b[92] = -32'sd64;
cb_b[93] = -32'sd62;
cb_b[94] = -32'sd60;
cb_b[95] = -32'sd58;
cb_b[96] = -32'sd57;
cb_b[97] = -32'sd55;
cb_b[98] = -32'sd53;
cb_b[99] = -32'sd51;
cb_b[100] = -32'sd50;
cb_b[101] = -32'sd48;
cb_b[102] = -32'sd46;
cb_b[103] = -32'sd44;
cb_b[104] = -32'sd43;
cb_b[105] = -32'sd41;
cb_b[106] = -32'sd39;
cb_b[107] = -32'sd37;
cb_b[108] = -32'sd35;
cb_b[109] = -32'sd34;
cb_b[110] = -32'sd32;
cb_b[111] = -32'sd30;
cb_b[112] = -32'sd28;
cb_b[113] = -32'sd27;
cb_b[114] = -32'sd25;
cb_b[115] = -32'sd23;
cb_b[116] = -32'sd21;
cb_b[117] = -32'sd19;
cb_b[118] = -32'sd18;
cb_b[119] = -32'sd16;
cb_b[120] = -32'sd14;
cb_b[121] = -32'sd12;
cb_b[122] = -32'sd11;
cb_b[123] = -32'sd9;
cb_b[124] = -32'sd7;
cb_b[125] = -32'sd5;
cb_b[126] = -32'sd4;
cb_b[127] = -32'sd2;
cb_b[128] = 32'sd0;
cb_b[129] = 32'sd2;
cb_b[130] = 32'sd4;
cb_b[131] = 32'sd5;
cb_b[132] = 32'sd7;
cb_b[133] = 32'sd9;
cb_b[134] = 32'sd11;
cb_b[135] = 32'sd12;
cb_b[136] = 32'sd14;
cb_b[137] = 32'sd16;
cb_b[138] = 32'sd18;
cb_b[139] = 32'sd19;
cb_b[140] = 32'sd21;
cb_b[141] = 32'sd23;
cb_b[142] = 32'sd25;
cb_b[143] = 32'sd27;
cb_b[144] = 32'sd28;
cb_b[145] = 32'sd30;
cb_b[146] = 32'sd32;
cb_b[147] = 32'sd34;
cb_b[148] = 32'sd35;
cb_b[149] = 32'sd37;
cb_b[150] = 32'sd39;
cb_b[151] = 32'sd41;
cb_b[152] = 32'sd43;
cb_b[153] = 32'sd44;
cb_b[154] = 32'sd46;
cb_b[155] = 32'sd48;
cb_b[156] = 32'sd50;
cb_b[157] = 32'sd51;
cb_b[158] = 32'sd53;
cb_b[159] = 32'sd55;
cb_b[160] = 32'sd57;
cb_b[161] = 32'sd58;
cb_b[162] = 32'sd60;
cb_b[163] = 32'sd62;
cb_b[164] = 32'sd64;
cb_b[165] = 32'sd66;
cb_b[166] = 32'sd67;
cb_b[167] = 32'sd69;
cb_b[168] = 32'sd71;
cb_b[169] = 32'sd73;
cb_b[170] = 32'sd74;
cb_b[171] = 32'sd76;
cb_b[172] = 32'sd78;
cb_b[173] = 32'sd80;
cb_b[174] = 32'sd82;
cb_b[175] = 32'sd83;
cb_b[176] = 32'sd85;
cb_b[177] = 32'sd87;
cb_b[178] = 32'sd89;
cb_b[179] = 32'sd90;
cb_b[180] = 32'sd92;
cb_b[181] = 32'sd94;
cb_b[182] = 32'sd96;
cb_b[183] = 32'sd97;
cb_b[184] = 32'sd99;
cb_b[185] = 32'sd101;
cb_b[186] = 32'sd103;
cb_b[187] = 32'sd105;
cb_b[188] = 32'sd106;
cb_b[189] = 32'sd108;
cb_b[190] = 32'sd110;
cb_b[191] = 32'sd112;
cb_b[192] = 32'sd113;
cb_b[193] = 32'sd115;
cb_b[194] = 32'sd117;
cb_b[195] = 32'sd119;
cb_b[196] = 32'sd120;
cb_b[197] = 32'sd122;
cb_b[198] = 32'sd124;
cb_b[199] = 32'sd126;
cb_b[200] = 32'sd128;
cb_b[201] = 32'sd129;
cb_b[202] = 32'sd131;
cb_b[203] = 32'sd133;
cb_b[204] = 32'sd135;
cb_b[205] = 32'sd136;
cb_b[206] = 32'sd138;
cb_b[207] = 32'sd140;
cb_b[208] = 32'sd142;
cb_b[209] = 32'sd144;
cb_b[210] = 32'sd145;
cb_b[211] = 32'sd147;
cb_b[212] = 32'sd149;
cb_b[213] = 32'sd151;
cb_b[214] = 32'sd152;
cb_b[215] = 32'sd154;
cb_b[216] = 32'sd156;
cb_b[217] = 32'sd158;
cb_b[218] = 32'sd159;
cb_b[219] = 32'sd161;
cb_b[220] = 32'sd163;
cb_b[221] = 32'sd165;
cb_b[222] = 32'sd167;
cb_b[223] = 32'sd168;
cb_b[224] = 32'sd170;
cb_b[225] = 32'sd172;
cb_b[226] = 32'sd174;
cb_b[227] = 32'sd175;
cb_b[228] = 32'sd177;
cb_b[229] = 32'sd179;
cb_b[230] = 32'sd181;
cb_b[231] = 32'sd183;
cb_b[232] = 32'sd184;
cb_b[233] = 32'sd186;
cb_b[234] = 32'sd188;
cb_b[235] = 32'sd190;
cb_b[236] = 32'sd191;
cb_b[237] = 32'sd193;
cb_b[238] = 32'sd195;
cb_b[239] = 32'sd197;
cb_b[240] = 32'sd198;
cb_b[241] = 32'sd200;
cb_b[242] = 32'sd202;
cb_b[243] = 32'sd204;
cb_b[244] = 32'sd206;
cb_b[245] = 32'sd207;
cb_b[246] = 32'sd209;
cb_b[247] = 32'sd211;
cb_b[248] = 32'sd213;
cb_b[249] = 32'sd214;
cb_b[250] = 32'sd216;
cb_b[251] = 32'sd218;
cb_b[252] = 32'sd220;
cb_b[253] = 32'sd222;
cb_b[254] = 32'sd223;
cb_b[255] = 32'sd225;

cb_g[0] = 32'sd2919680;
cb_g[1] = 32'sd2897126;
cb_g[2] = 32'sd2874572;
cb_g[3] = 32'sd2852018;
cb_g[4] = 32'sd2829464;
cb_g[5] = 32'sd2806910;
cb_g[6] = 32'sd2784356;
cb_g[7] = 32'sd2761802;
cb_g[8] = 32'sd2739248;
cb_g[9] = 32'sd2716694;
cb_g[10] = 32'sd2694140;
cb_g[11] = 32'sd2671586;
cb_g[12] = 32'sd2649032;
cb_g[13] = 32'sd2626478;
cb_g[14] = 32'sd2603924;
cb_g[15] = 32'sd2581370;
cb_g[16] = 32'sd2558816;
cb_g[17] = 32'sd2536262;
cb_g[18] = 32'sd2513708;
cb_g[19] = 32'sd2491154;
cb_g[20] = 32'sd2468600;
cb_g[21] = 32'sd2446046;
cb_g[22] = 32'sd2423492;
cb_g[23] = 32'sd2400938;
cb_g[24] = 32'sd2378384;
cb_g[25] = 32'sd2355830;
cb_g[26] = 32'sd2333276;
cb_g[27] = 32'sd2310722;
cb_g[28] = 32'sd2288168;
cb_g[29] = 32'sd2265614;
cb_g[30] = 32'sd2243060;
cb_g[31] = 32'sd2220506;
cb_g[32] = 32'sd2197952;
cb_g[33] = 32'sd2175398;
cb_g[34] = 32'sd2152844;
cb_g[35] = 32'sd2130290;
cb_g[36] = 32'sd2107736;
cb_g[37] = 32'sd2085182;
cb_g[38] = 32'sd2062628;
cb_g[39] = 32'sd2040074;
cb_g[40] = 32'sd2017520;
cb_g[41] = 32'sd1994966;
cb_g[42] = 32'sd1972412;
cb_g[43] = 32'sd1949858;
cb_g[44] = 32'sd1927304;
cb_g[45] = 32'sd1904750;
cb_g[46] = 32'sd1882196;
cb_g[47] = 32'sd1859642;
cb_g[48] = 32'sd1837088;
cb_g[49] = 32'sd1814534;
cb_g[50] = 32'sd1791980;
cb_g[51] = 32'sd1769426;
cb_g[52] = 32'sd1746872;
cb_g[53] = 32'sd1724318;
cb_g[54] = 32'sd1701764;
cb_g[55] = 32'sd1679210;
cb_g[56] = 32'sd1656656;
cb_g[57] = 32'sd1634102;
cb_g[58] = 32'sd1611548;
cb_g[59] = 32'sd1588994;
cb_g[60] = 32'sd1566440;
cb_g[61] = 32'sd1543886;
cb_g[62] = 32'sd1521332;
cb_g[63] = 32'sd1498778;
cb_g[64] = 32'sd1476224;
cb_g[65] = 32'sd1453670;
cb_g[66] = 32'sd1431116;
cb_g[67] = 32'sd1408562;
cb_g[68] = 32'sd1386008;
cb_g[69] = 32'sd1363454;
cb_g[70] = 32'sd1340900;
cb_g[71] = 32'sd1318346;
cb_g[72] = 32'sd1295792;
cb_g[73] = 32'sd1273238;
cb_g[74] = 32'sd1250684;
cb_g[75] = 32'sd1228130;
cb_g[76] = 32'sd1205576;
cb_g[77] = 32'sd1183022;
cb_g[78] = 32'sd1160468;
cb_g[79] = 32'sd1137914;
cb_g[80] = 32'sd1115360;
cb_g[81] = 32'sd1092806;
cb_g[82] = 32'sd1070252;
cb_g[83] = 32'sd1047698;
cb_g[84] = 32'sd1025144;
cb_g[85] = 32'sd1002590;
cb_g[86] = 32'sd980036;
cb_g[87] = 32'sd957482;
cb_g[88] = 32'sd934928;
cb_g[89] = 32'sd912374;
cb_g[90] = 32'sd889820;
cb_g[91] = 32'sd867266;
cb_g[92] = 32'sd844712;
cb_g[93] = 32'sd822158;
cb_g[94] = 32'sd799604;
cb_g[95] = 32'sd777050;
cb_g[96] = 32'sd754496;
cb_g[97] = 32'sd731942;
cb_g[98] = 32'sd709388;
cb_g[99] = 32'sd686834;
cb_g[100] = 32'sd664280;
cb_g[101] = 32'sd641726;
cb_g[102] = 32'sd619172;
cb_g[103] = 32'sd596618;
cb_g[104] = 32'sd574064;
cb_g[105] = 32'sd551510;
cb_g[106] = 32'sd528956;
cb_g[107] = 32'sd506402;
cb_g[108] = 32'sd483848;
cb_g[109] = 32'sd461294;
cb_g[110] = 32'sd438740;
cb_g[111] = 32'sd416186;
cb_g[112] = 32'sd393632;
cb_g[113] = 32'sd371078;
cb_g[114] = 32'sd348524;
cb_g[115] = 32'sd325970;
cb_g[116] = 32'sd303416;
cb_g[117] = 32'sd280862;
cb_g[118] = 32'sd258308;
cb_g[119] = 32'sd235754;
cb_g[120] = 32'sd213200;
cb_g[121] = 32'sd190646;
cb_g[122] = 32'sd168092;
cb_g[123] = 32'sd145538;
cb_g[124] = 32'sd122984;
cb_g[125] = 32'sd100430;
cb_g[126] = 32'sd77876;
cb_g[127] = 32'sd55322;
cb_g[128] = 32'sd32768;
cb_g[129] = 32'sd10214;
cb_g[130] = -32'sd12340;
cb_g[131] = -32'sd34894;
cb_g[132] = -32'sd57448;
cb_g[133] = -32'sd80002;
cb_g[134] = -32'sd102556;
cb_g[135] = -32'sd125110;
cb_g[136] = -32'sd147664;
cb_g[137] = -32'sd170218;
cb_g[138] = -32'sd192772;
cb_g[139] = -32'sd215326;
cb_g[140] = -32'sd237880;
cb_g[141] = -32'sd260434;
cb_g[142] = -32'sd282988;
cb_g[143] = -32'sd305542;
cb_g[144] = -32'sd328096;
cb_g[145] = -32'sd350650;
cb_g[146] = -32'sd373204;
cb_g[147] = -32'sd395758;
cb_g[148] = -32'sd418312;
cb_g[149] = -32'sd440866;
cb_g[150] = -32'sd463420;
cb_g[151] = -32'sd485974;
cb_g[152] = -32'sd508528;
cb_g[153] = -32'sd531082;
cb_g[154] = -32'sd553636;
cb_g[155] = -32'sd576190;
cb_g[156] = -32'sd598744;
cb_g[157] = -32'sd621298;
cb_g[158] = -32'sd643852;
cb_g[159] = -32'sd666406;
cb_g[160] = -32'sd688960;
cb_g[161] = -32'sd711514;
cb_g[162] = -32'sd734068;
cb_g[163] = -32'sd756622;
cb_g[164] = -32'sd779176;
cb_g[165] = -32'sd801730;
cb_g[166] = -32'sd824284;
cb_g[167] = -32'sd846838;
cb_g[168] = -32'sd869392;
cb_g[169] = -32'sd891946;
cb_g[170] = -32'sd914500;
cb_g[171] = -32'sd937054;
cb_g[172] = -32'sd959608;
cb_g[173] = -32'sd982162;
cb_g[174] = -32'sd1004716;
cb_g[175] = -32'sd1027270;
cb_g[176] = -32'sd1049824;
cb_g[177] = -32'sd1072378;
cb_g[178] = -32'sd1094932;
cb_g[179] = -32'sd1117486;
cb_g[180] = -32'sd1140040;
cb_g[181] = -32'sd1162594;
cb_g[182] = -32'sd1185148;
cb_g[183] = -32'sd1207702;
cb_g[184] = -32'sd1230256;
cb_g[185] = -32'sd1252810;
cb_g[186] = -32'sd1275364;
cb_g[187] = -32'sd1297918;
cb_g[188] = -32'sd1320472;
cb_g[189] = -32'sd1343026;
cb_g[190] = -32'sd1365580;
cb_g[191] = -32'sd1388134;
cb_g[192] = -32'sd1410688;
cb_g[193] = -32'sd1433242;
cb_g[194] = -32'sd1455796;
cb_g[195] = -32'sd1478350;
cb_g[196] = -32'sd1500904;
cb_g[197] = -32'sd1523458;
cb_g[198] = -32'sd1546012;
cb_g[199] = -32'sd1568566;
cb_g[200] = -32'sd1591120;
cb_g[201] = -32'sd1613674;
cb_g[202] = -32'sd1636228;
cb_g[203] = -32'sd1658782;
cb_g[204] = -32'sd1681336;
cb_g[205] = -32'sd1703890;
cb_g[206] = -32'sd1726444;
cb_g[207] = -32'sd1748998;
cb_g[208] = -32'sd1771552;
cb_g[209] = -32'sd1794106;
cb_g[210] = -32'sd1816660;
cb_g[211] = -32'sd1839214;
cb_g[212] = -32'sd1861768;
cb_g[213] = -32'sd1884322;
cb_g[214] = -32'sd1906876;
cb_g[215] = -32'sd1929430;
cb_g[216] = -32'sd1951984;
cb_g[217] = -32'sd1974538;
cb_g[218] = -32'sd1997092;
cb_g[219] = -32'sd2019646;
cb_g[220] = -32'sd2042200;
cb_g[221] = -32'sd2064754;
cb_g[222] = -32'sd2087308;
cb_g[223] = -32'sd2109862;
cb_g[224] = -32'sd2132416;
cb_g[225] = -32'sd2154970;
cb_g[226] = -32'sd2177524;
cb_g[227] = -32'sd2200078;
cb_g[228] = -32'sd2222632;
cb_g[229] = -32'sd2245186;
cb_g[230] = -32'sd2267740;
cb_g[231] = -32'sd2290294;
cb_g[232] = -32'sd2312848;
cb_g[233] = -32'sd2335402;
cb_g[234] = -32'sd2357956;
cb_g[235] = -32'sd2380510;
cb_g[236] = -32'sd2403064;
cb_g[237] = -32'sd2425618;
cb_g[238] = -32'sd2448172;
cb_g[239] = -32'sd2470726;
cb_g[240] = -32'sd2493280;
cb_g[241] = -32'sd2515834;
cb_g[242] = -32'sd2538388;
cb_g[243] = -32'sd2560942;
cb_g[244] = -32'sd2583496;
cb_g[245] = -32'sd2606050;
cb_g[246] = -32'sd2628604;
cb_g[247] = -32'sd2651158;
cb_g[248] = -32'sd2673712;
cb_g[249] = -32'sd2696266;
cb_g[250] = -32'sd2718820;
cb_g[251] = -32'sd2741374;
cb_g[252] = -32'sd2763928;
cb_g[253] = -32'sd2786482;
cb_g[254] = -32'sd2809036;
cb_g[255] = -32'sd2831590;



end

always 
begin

dataa_reg = dataa;
datab_reg = datab;

y = dataa_reg[7:0];
cr = datab_reg[7:0];
cb = datab_reg[15:8];

R = y + cr_r[cr];
G = y + ((cb_g[cb] + cr_g[cr]) >> 16);
B = y + cb_b[cb];

result = {R,G,B}; 
end
endmodule

